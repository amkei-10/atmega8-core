/home/mario/Dropbox/ProzessorDesign/progmem_hex2vhd/pkg_instrmem.vhd