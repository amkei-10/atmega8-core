library ieee;
use ieee.std_logic_1164.all;
-- ---------------------------------------------------------------------------------
-- Memory initialisation package
-- ---------------------------------------------------------------------------------
package pkg_instrmem is

	type t_instrMem   is array(0 to 512-1) of std_logic_vector(15 downto 0);
	constant PROGMEM : t_instrMem := (
		"1110000001100100",
		"0010011111111111",
		"1110001111100011",
		"1000000010110000",
		"1110001111100110",
		"1000000010100000",
		"1110001111100101",
		"1000001010110000",
		"1101000001001110",
		"1110001111101000",
		"1000001010100000",
		"0010110100011010",
		"0111000000011111",
		"1101000000011111",
		"1110010011100001",
		"1000001100000000",
		"0010110100011010",
		"1001010100010110",
		"1001010100010110",
		"1001010100010110",
		"1001010100010110",
		"1101000000010111",
		"1110010011100010",
		"1000001100000000",
		"0010110100011011",
		"0111000000011111",
		"1101000000010010",
		"1110010011100011",
		"1000001100000000",
		"0010110100011011",
		"1001010100010110",
		"1001010100010110",
		"1001010100010110",
		"1001010100010110",
		"1101000000001010",
		"1110010011100100",
		"1000001100000000",
		"1110010011100000",
		"0011000101100000",
		"1111010000001001",
		"1110000001100001",
		"1000001101100000",
		"0000111101100110",
		"1101000000101011",
		"1100111111010100",
		"0011000000010000",
		"1111010000010001",
		"1110001100001111",
		"1001010100001000",
		"0011000000010001",
		"1111010000010001",
		"1110000000000110",
		"1001010100001000",
		"0011000000010010",
		"1111010000010001",
		"1110010100001011",
		"1001010100001000",
		"0011000000010011",
		"1111010000010001",
		"1110010000001111",
		"1001010100001000",
		"0011000000010100",
		"1111010000010001",
		"1110011000000110",
		"1001010100001000",
		"0011000000010101",
		"1111010000010001",
		"1110011000001101",
		"1001010100001000",
		"0011000000010110",
		"1111010000010001",
		"1110011100001101",
		"1001010100001000",
		"0011000000010111",
		"1111010000010001",
		"1110000000000111",
		"1001010100001000",
		"0011000000011000",
		"1111010000010001",
		"1110011100001111",
		"1001010100001000",
		"0011000000011001",
		"1111010000010001",
		"1110011000001111",
		"1001010100001000",
		"1110111100001001",
		"1001010100001000",
		"0010011100100010",
		"0010011100110011",
		"0010011101000100",
		"1001010101001010",
		"1111011111110001",
		"1001010100111010",
		"1111011111011001",
		"1001010100101010",
		"1111011111000001",
		"1001010100001000",
		
		others => (others => '0')
	);

end package pkg_instrmem;
